* parameter sweep
* code obtained from ngspice sourceforge forum user marcel hendrix
* extra comment

* this works when this is the CURRENT ...thing
* have to restart ngspice
* resistive divider , R1 swept from start_r to stop_r
VDD 1 0 DC=1V
R1  1 2 1k
R2  2 0 1k

.control
let start_r = 1k
let stop_r  = 10k
let delta_r = 1k
let r_act   = start_r
* loop
echo parameter sweep > result.txt
while r_act le stop_r
  alter r1 r_act
  op
  *let expect = 1k/(r_act+1k)
  *echo $&r_act $&v(2) $&expect >> result.txt
  print v(2)
  let r_act = r_act + delta_r
end
.endc

.end
