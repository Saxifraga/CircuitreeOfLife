* High pass filter
.ac dec 10 1 1e5
.control
save all
run
write
.endc

V1 1 0 ac 1
C1 1 2 0.0952335570127u
R2 2 0 0.495327116872k
C3 2 3 0.878964408256u
C4 3 0 0.884476082001u
.END